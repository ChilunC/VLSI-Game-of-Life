magic
tech scmos
timestamp 1519843622
<< m2contact >>
rect -2 -2 2 2
<< end >>
