magic
tech scmos
timestamp 1519843622
<< nwell >>
rect -8 48 32 105
<< ntransistor >>
rect 7 6 9 26
rect 12 6 14 26
<< ptransistor >>
rect 7 74 9 94
rect 15 74 17 94
<< ndiffusion >>
rect 2 25 7 26
rect 6 6 7 25
rect 9 6 12 26
rect 14 25 19 26
rect 14 6 15 25
<< pdiffusion >>
rect 2 93 7 94
rect 6 74 7 93
rect 9 93 15 94
rect 9 74 10 93
rect 14 74 15 93
rect 17 93 22 94
rect 17 74 18 93
<< ndcontact >>
rect 2 6 6 25
rect 15 6 19 25
<< pdcontact >>
rect 2 74 6 93
rect 10 74 14 93
rect 18 74 22 93
<< psubstratepcontact >>
rect -2 -2 2 2
rect 14 -2 18 2
<< nsubstratencontact >>
rect -2 98 2 102
rect 14 98 18 102
<< polysilicon >>
rect 7 94 9 96
rect 15 94 17 96
rect 7 33 9 74
rect 6 29 9 33
rect 15 61 17 74
rect 15 57 18 61
rect 15 29 17 57
rect 7 26 9 29
rect 12 27 17 29
rect 12 26 14 27
rect 7 4 9 6
rect 12 4 14 6
<< polycontact >>
rect 2 29 6 33
rect 18 57 22 61
<< metal1 >>
rect -2 102 26 103
rect 2 98 14 102
rect 18 98 26 102
rect -2 97 26 98
rect 2 93 6 97
rect 10 93 14 94
rect 18 93 22 97
rect 2 33 6 37
rect 10 26 14 74
rect 18 53 22 57
rect 2 25 6 26
rect 10 25 19 26
rect 10 23 15 25
rect 2 3 6 6
rect -2 2 26 3
rect 2 -2 14 2
rect 18 -2 26 2
rect -2 -3 26 -2
<< m1p >>
rect 18 53 22 57
rect 10 43 14 47
rect 2 33 6 37
<< labels >>
rlabel metal1 4 100 4 100 4 vdd
rlabel metal1 12 45 12 45 4 Y
rlabel metal1 4 0 4 0 4 gnd
rlabel metal1 4 35 4 35 4 A
rlabel metal1 20 55 20 55 4 B
<< end >>
